module case_top
  (
   input clk,
   input [8:0] neighbors,
   output result
   );
  

  reg [8:0]   neighbors_r;
  reg	      wdata;
  assign result = wdata;
  
  always @ (posedge clk) begin
    neighbors_r <= neighbors;
  end

  always @(posedge clk) begin
    case(neighbors_r)
      9'b000_000_000: wdata <= 1'b0;
      9'b000_000_001: wdata <= 1'b0;
      9'b000_000_010: wdata <= 1'b0;
      9'b000_000_011: wdata <= 1'b0;
      9'b000_000_100: wdata <= 1'b0;
      9'b000_000_101: wdata <= 1'b0;
      9'b000_000_110: wdata <= 1'b0;
      9'b000_000_111: wdata <= 1'b1;
      9'b000_001_000: wdata <= 1'b0;
      9'b000_001_001: wdata <= 1'b0;
      9'b000_001_010: wdata <= 1'b0;
      9'b000_001_011: wdata <= 1'b1;
      9'b000_001_100: wdata <= 1'b0;
      9'b000_001_101: wdata <= 1'b1;
      9'b000_001_110: wdata <= 1'b1;
      9'b000_001_111: wdata <= 1'b0;
      9'b000_010_000: wdata <= 1'b0;
      9'b000_010_001: wdata <= 1'b0;
      9'b000_010_010: wdata <= 1'b0;
      9'b000_010_011: wdata <= 1'b1;
      9'b000_010_100: wdata <= 1'b0;
      9'b000_010_101: wdata <= 1'b1;
      9'b000_010_110: wdata <= 1'b1;
      9'b000_010_111: wdata <= 1'b1;
      9'b000_011_000: wdata <= 1'b0;
      9'b000_011_001: wdata <= 1'b1;
      9'b000_011_010: wdata <= 1'b1;
      9'b000_011_011: wdata <= 1'b1;
      9'b000_011_100: wdata <= 1'b1;
      9'b000_011_101: wdata <= 1'b1;
      9'b000_011_110: wdata <= 1'b1;
      9'b000_011_111: wdata <= 1'b0;
      9'b000_100_000: wdata <= 1'b0;
      9'b000_100_001: wdata <= 1'b0;
      9'b000_100_010: wdata <= 1'b0;
      9'b000_100_011: wdata <= 1'b1;
      9'b000_100_100: wdata <= 1'b0;
      9'b000_100_101: wdata <= 1'b1;
      9'b000_100_110: wdata <= 1'b1;
      9'b000_100_111: wdata <= 1'b0;
      9'b000_101_000: wdata <= 1'b0;
      9'b000_101_001: wdata <= 1'b1;
      9'b000_101_010: wdata <= 1'b1;
      9'b000_101_011: wdata <= 1'b0;
      9'b000_101_100: wdata <= 1'b1;
      9'b000_101_101: wdata <= 1'b0;
      9'b000_101_110: wdata <= 1'b0;
      9'b000_101_111: wdata <= 1'b0;
      9'b000_110_000: wdata <= 1'b0;
      9'b000_110_001: wdata <= 1'b1;
      9'b000_110_010: wdata <= 1'b1;
      9'b000_110_011: wdata <= 1'b1;
      9'b000_110_100: wdata <= 1'b1;
      9'b000_110_101: wdata <= 1'b1;
      9'b000_110_110: wdata <= 1'b1;
      9'b000_110_111: wdata <= 1'b0;
      9'b000_111_000: wdata <= 1'b1;
      9'b000_111_001: wdata <= 1'b1;
      9'b000_111_010: wdata <= 1'b1;
      9'b000_111_011: wdata <= 1'b0;
      9'b000_111_100: wdata <= 1'b1;
      9'b000_111_101: wdata <= 1'b0;
      9'b000_111_110: wdata <= 1'b0;
      9'b000_111_111: wdata <= 1'b0;
      9'b001_000_000: wdata <= 1'b0;
      9'b001_000_001: wdata <= 1'b0;
      9'b001_000_010: wdata <= 1'b0;
      9'b001_000_011: wdata <= 1'b1;
      9'b001_000_100: wdata <= 1'b0;
      9'b001_000_101: wdata <= 1'b1;
      9'b001_000_110: wdata <= 1'b1;
      9'b001_000_111: wdata <= 1'b0;
      9'b001_001_000: wdata <= 1'b0;
      9'b001_001_001: wdata <= 1'b1;
      9'b001_001_010: wdata <= 1'b1;
      9'b001_001_011: wdata <= 1'b0;
      9'b001_001_100: wdata <= 1'b1;
      9'b001_001_101: wdata <= 1'b0;
      9'b001_001_110: wdata <= 1'b0;
      9'b001_001_111: wdata <= 1'b0;
      9'b001_010_000: wdata <= 1'b0;
      9'b001_010_001: wdata <= 1'b1;
      9'b001_010_010: wdata <= 1'b1;
      9'b001_010_011: wdata <= 1'b1;
      9'b001_010_100: wdata <= 1'b1;
      9'b001_010_101: wdata <= 1'b1;
      9'b001_010_110: wdata <= 1'b1;
      9'b001_010_111: wdata <= 1'b0;
      9'b001_011_000: wdata <= 1'b1;
      9'b001_011_001: wdata <= 1'b1;
      9'b001_011_010: wdata <= 1'b1;
      9'b001_011_011: wdata <= 1'b0;
      9'b001_011_100: wdata <= 1'b1;
      9'b001_011_101: wdata <= 1'b0;
      9'b001_011_110: wdata <= 1'b0;
      9'b001_011_111: wdata <= 1'b0;
      9'b001_100_000: wdata <= 1'b0;
      9'b001_100_001: wdata <= 1'b1;
      9'b001_100_010: wdata <= 1'b1;
      9'b001_100_011: wdata <= 1'b0;
      9'b001_100_100: wdata <= 1'b1;
      9'b001_100_101: wdata <= 1'b0;
      9'b001_100_110: wdata <= 1'b0;
      9'b001_100_111: wdata <= 1'b0;
      9'b001_101_000: wdata <= 1'b1;
      9'b001_101_001: wdata <= 1'b0;
      9'b001_101_010: wdata <= 1'b0;
      9'b001_101_011: wdata <= 1'b0;
      9'b001_101_100: wdata <= 1'b0;
      9'b001_101_101: wdata <= 1'b0;
      9'b001_101_110: wdata <= 1'b0;
      9'b001_101_111: wdata <= 1'b0;
      9'b001_110_000: wdata <= 1'b1;
      9'b001_110_001: wdata <= 1'b1;
      9'b001_110_010: wdata <= 1'b1;
      9'b001_110_011: wdata <= 1'b0;
      9'b001_110_100: wdata <= 1'b1;
      9'b001_110_101: wdata <= 1'b0;
      9'b001_110_110: wdata <= 1'b0;
      9'b001_110_111: wdata <= 1'b0;
      9'b001_111_000: wdata <= 1'b1;
      9'b001_111_001: wdata <= 1'b0;
      9'b001_111_010: wdata <= 1'b0;
      9'b001_111_011: wdata <= 1'b0;
      9'b001_111_100: wdata <= 1'b0;
      9'b001_111_101: wdata <= 1'b0;
      9'b001_111_110: wdata <= 1'b0;
      9'b001_111_111: wdata <= 1'b0;
      9'b010_000_000: wdata <= 1'b0;
      9'b010_000_001: wdata <= 1'b0;
      9'b010_000_010: wdata <= 1'b0;
      9'b010_000_011: wdata <= 1'b1;
      9'b010_000_100: wdata <= 1'b0;
      9'b010_000_101: wdata <= 1'b1;
      9'b010_000_110: wdata <= 1'b1;
      9'b010_000_111: wdata <= 1'b0;
      9'b010_001_000: wdata <= 1'b0;
      9'b010_001_001: wdata <= 1'b1;
      9'b010_001_010: wdata <= 1'b1;
      9'b010_001_011: wdata <= 1'b0;
      9'b010_001_100: wdata <= 1'b1;
      9'b010_001_101: wdata <= 1'b0;
      9'b010_001_110: wdata <= 1'b0;
      9'b010_001_111: wdata <= 1'b0;
      9'b010_010_000: wdata <= 1'b0;
      9'b010_010_001: wdata <= 1'b1;
      9'b010_010_010: wdata <= 1'b1;
      9'b010_010_011: wdata <= 1'b1;
      9'b010_010_100: wdata <= 1'b1;
      9'b010_010_101: wdata <= 1'b1;
      9'b010_010_110: wdata <= 1'b1;
      9'b010_010_111: wdata <= 1'b0;
      9'b010_011_000: wdata <= 1'b1;
      9'b010_011_001: wdata <= 1'b1;
      9'b010_011_010: wdata <= 1'b1;
      9'b010_011_011: wdata <= 1'b0;
      9'b010_011_100: wdata <= 1'b1;
      9'b010_011_101: wdata <= 1'b0;
      9'b010_011_110: wdata <= 1'b0;
      9'b010_011_111: wdata <= 1'b0;
      9'b010_100_000: wdata <= 1'b0;
      9'b010_100_001: wdata <= 1'b1;
      9'b010_100_010: wdata <= 1'b1;
      9'b010_100_011: wdata <= 1'b0;
      9'b010_100_100: wdata <= 1'b1;
      9'b010_100_101: wdata <= 1'b0;
      9'b010_100_110: wdata <= 1'b0;
      9'b010_100_111: wdata <= 1'b0;
      9'b010_101_000: wdata <= 1'b1;
      9'b010_101_001: wdata <= 1'b0;
      9'b010_101_010: wdata <= 1'b0;
      9'b010_101_011: wdata <= 1'b0;
      9'b010_101_100: wdata <= 1'b0;
      9'b010_101_101: wdata <= 1'b0;
      9'b010_101_110: wdata <= 1'b0;
      9'b010_101_111: wdata <= 1'b0;
      9'b010_110_000: wdata <= 1'b1;
      9'b010_110_001: wdata <= 1'b1;
      9'b010_110_010: wdata <= 1'b1;
      9'b010_110_011: wdata <= 1'b0;
      9'b010_110_100: wdata <= 1'b1;
      9'b010_110_101: wdata <= 1'b0;
      9'b010_110_110: wdata <= 1'b0;
      9'b010_110_111: wdata <= 1'b0;
      9'b010_111_000: wdata <= 1'b1;
      9'b010_111_001: wdata <= 1'b0;
      9'b010_111_010: wdata <= 1'b0;
      9'b010_111_011: wdata <= 1'b0;
      9'b010_111_100: wdata <= 1'b0;
      9'b010_111_101: wdata <= 1'b0;
      9'b010_111_110: wdata <= 1'b0;
      9'b010_111_111: wdata <= 1'b0;
      9'b011_000_000: wdata <= 1'b0;
      9'b011_000_001: wdata <= 1'b1;
      9'b011_000_010: wdata <= 1'b1;
      9'b011_000_011: wdata <= 1'b0;
      9'b011_000_100: wdata <= 1'b1;
      9'b011_000_101: wdata <= 1'b0;
      9'b011_000_110: wdata <= 1'b0;
      9'b011_000_111: wdata <= 1'b0;
      9'b011_001_000: wdata <= 1'b1;
      9'b011_001_001: wdata <= 1'b0;
      9'b011_001_010: wdata <= 1'b0;
      9'b011_001_011: wdata <= 1'b0;
      9'b011_001_100: wdata <= 1'b0;
      9'b011_001_101: wdata <= 1'b0;
      9'b011_001_110: wdata <= 1'b0;
      9'b011_001_111: wdata <= 1'b0;
      9'b011_010_000: wdata <= 1'b1;
      9'b011_010_001: wdata <= 1'b1;
      9'b011_010_010: wdata <= 1'b1;
      9'b011_010_011: wdata <= 1'b0;
      9'b011_010_100: wdata <= 1'b1;
      9'b011_010_101: wdata <= 1'b0;
      9'b011_010_110: wdata <= 1'b0;
      9'b011_010_111: wdata <= 1'b0;
      9'b011_011_000: wdata <= 1'b1;
      9'b011_011_001: wdata <= 1'b0;
      9'b011_011_010: wdata <= 1'b0;
      9'b011_011_011: wdata <= 1'b0;
      9'b011_011_100: wdata <= 1'b0;
      9'b011_011_101: wdata <= 1'b0;
      9'b011_011_110: wdata <= 1'b0;
      9'b011_011_111: wdata <= 1'b0;
      9'b011_100_000: wdata <= 1'b1;
      9'b011_100_001: wdata <= 1'b0;
      9'b011_100_010: wdata <= 1'b0;
      9'b011_100_011: wdata <= 1'b0;
      9'b011_100_100: wdata <= 1'b0;
      9'b011_100_101: wdata <= 1'b0;
      9'b011_100_110: wdata <= 1'b0;
      9'b011_100_111: wdata <= 1'b0;
      9'b011_101_000: wdata <= 1'b0;
      9'b011_101_001: wdata <= 1'b0;
      9'b011_101_010: wdata <= 1'b0;
      9'b011_101_011: wdata <= 1'b0;
      9'b011_101_100: wdata <= 1'b0;
      9'b011_101_101: wdata <= 1'b0;
      9'b011_101_110: wdata <= 1'b0;
      9'b011_101_111: wdata <= 1'b0;
      9'b011_110_000: wdata <= 1'b1;
      9'b011_110_001: wdata <= 1'b0;
      9'b011_110_010: wdata <= 1'b0;
      9'b011_110_011: wdata <= 1'b0;
      9'b011_110_100: wdata <= 1'b0;
      9'b011_110_101: wdata <= 1'b0;
      9'b011_110_110: wdata <= 1'b0;
      9'b011_110_111: wdata <= 1'b0;
      9'b011_111_000: wdata <= 1'b0;
      9'b011_111_001: wdata <= 1'b0;
      9'b011_111_010: wdata <= 1'b0;
      9'b011_111_011: wdata <= 1'b0;
      9'b011_111_100: wdata <= 1'b0;
      9'b011_111_101: wdata <= 1'b0;
      9'b011_111_110: wdata <= 1'b0;
      9'b011_111_111: wdata <= 1'b0;
      9'b100_000_000: wdata <= 1'b0;
      9'b100_000_001: wdata <= 1'b0;
      9'b100_000_010: wdata <= 1'b0;
      9'b100_000_011: wdata <= 1'b1;
      9'b100_000_100: wdata <= 1'b0;
      9'b100_000_101: wdata <= 1'b1;
      9'b100_000_110: wdata <= 1'b1;
      9'b100_000_111: wdata <= 1'b0;
      9'b100_001_000: wdata <= 1'b0;
      9'b100_001_001: wdata <= 1'b1;
      9'b100_001_010: wdata <= 1'b1;
      9'b100_001_011: wdata <= 1'b0;
      9'b100_001_100: wdata <= 1'b1;
      9'b100_001_101: wdata <= 1'b0;
      9'b100_001_110: wdata <= 1'b0;
      9'b100_001_111: wdata <= 1'b0;
      9'b100_010_000: wdata <= 1'b0;
      9'b100_010_001: wdata <= 1'b1;
      9'b100_010_010: wdata <= 1'b1;
      9'b100_010_011: wdata <= 1'b1;
      9'b100_010_100: wdata <= 1'b1;
      9'b100_010_101: wdata <= 1'b1;
      9'b100_010_110: wdata <= 1'b1;
      9'b100_010_111: wdata <= 1'b0;
      9'b100_011_000: wdata <= 1'b1;
      9'b100_011_001: wdata <= 1'b1;
      9'b100_011_010: wdata <= 1'b1;
      9'b100_011_011: wdata <= 1'b0;
      9'b100_011_100: wdata <= 1'b1;
      9'b100_011_101: wdata <= 1'b0;
      9'b100_011_110: wdata <= 1'b0;
      9'b100_011_111: wdata <= 1'b0;
      9'b100_100_000: wdata <= 1'b0;
      9'b100_100_001: wdata <= 1'b1;
      9'b100_100_010: wdata <= 1'b1;
      9'b100_100_011: wdata <= 1'b0;
      9'b100_100_100: wdata <= 1'b1;
      9'b100_100_101: wdata <= 1'b0;
      9'b100_100_110: wdata <= 1'b0;
      9'b100_100_111: wdata <= 1'b0;
      9'b100_101_000: wdata <= 1'b1;
      9'b100_101_001: wdata <= 1'b0;
      9'b100_101_010: wdata <= 1'b0;
      9'b100_101_011: wdata <= 1'b0;
      9'b100_101_100: wdata <= 1'b0;
      9'b100_101_101: wdata <= 1'b0;
      9'b100_101_110: wdata <= 1'b0;
      9'b100_101_111: wdata <= 1'b0;
      9'b100_110_000: wdata <= 1'b1;
      9'b100_110_001: wdata <= 1'b1;
      9'b100_110_010: wdata <= 1'b1;
      9'b100_110_011: wdata <= 1'b0;
      9'b100_110_100: wdata <= 1'b1;
      9'b100_110_101: wdata <= 1'b0;
      9'b100_110_110: wdata <= 1'b0;
      9'b100_110_111: wdata <= 1'b0;
      9'b100_111_000: wdata <= 1'b1;
      9'b100_111_001: wdata <= 1'b0;
      9'b100_111_010: wdata <= 1'b0;
      9'b100_111_011: wdata <= 1'b0;
      9'b100_111_100: wdata <= 1'b0;
      9'b100_111_101: wdata <= 1'b0;
      9'b100_111_110: wdata <= 1'b0;
      9'b100_111_111: wdata <= 1'b0;
      9'b101_000_000: wdata <= 1'b0;
      9'b101_000_001: wdata <= 1'b1;
      9'b101_000_010: wdata <= 1'b1;
      9'b101_000_011: wdata <= 1'b0;
      9'b101_000_100: wdata <= 1'b1;
      9'b101_000_101: wdata <= 1'b0;
      9'b101_000_110: wdata <= 1'b0;
      9'b101_000_111: wdata <= 1'b0;
      9'b101_001_000: wdata <= 1'b1;
      9'b101_001_001: wdata <= 1'b0;
      9'b101_001_010: wdata <= 1'b0;
      9'b101_001_011: wdata <= 1'b0;
      9'b101_001_100: wdata <= 1'b0;
      9'b101_001_101: wdata <= 1'b0;
      9'b101_001_110: wdata <= 1'b0;
      9'b101_001_111: wdata <= 1'b0;
      9'b101_010_000: wdata <= 1'b1;
      9'b101_010_001: wdata <= 1'b1;
      9'b101_010_010: wdata <= 1'b1;
      9'b101_010_011: wdata <= 1'b0;
      9'b101_010_100: wdata <= 1'b1;
      9'b101_010_101: wdata <= 1'b0;
      9'b101_010_110: wdata <= 1'b0;
      9'b101_010_111: wdata <= 1'b0;
      9'b101_011_000: wdata <= 1'b1;
      9'b101_011_001: wdata <= 1'b0;
      9'b101_011_010: wdata <= 1'b0;
      9'b101_011_011: wdata <= 1'b0;
      9'b101_011_100: wdata <= 1'b0;
      9'b101_011_101: wdata <= 1'b0;
      9'b101_011_110: wdata <= 1'b0;
      9'b101_011_111: wdata <= 1'b0;
      9'b101_100_000: wdata <= 1'b1;
      9'b101_100_001: wdata <= 1'b0;
      9'b101_100_010: wdata <= 1'b0;
      9'b101_100_011: wdata <= 1'b0;
      9'b101_100_100: wdata <= 1'b0;
      9'b101_100_101: wdata <= 1'b0;
      9'b101_100_110: wdata <= 1'b0;
      9'b101_100_111: wdata <= 1'b0;
      9'b101_101_000: wdata <= 1'b0;
      9'b101_101_001: wdata <= 1'b0;
      9'b101_101_010: wdata <= 1'b0;
      9'b101_101_011: wdata <= 1'b0;
      9'b101_101_100: wdata <= 1'b0;
      9'b101_101_101: wdata <= 1'b0;
      9'b101_101_110: wdata <= 1'b0;
      9'b101_101_111: wdata <= 1'b0;
      9'b101_110_000: wdata <= 1'b1;
      9'b101_110_001: wdata <= 1'b0;
      9'b101_110_010: wdata <= 1'b0;
      9'b101_110_011: wdata <= 1'b0;
      9'b101_110_100: wdata <= 1'b0;
      9'b101_110_101: wdata <= 1'b0;
      9'b101_110_110: wdata <= 1'b0;
      9'b101_110_111: wdata <= 1'b0;
      9'b101_111_000: wdata <= 1'b0;
      9'b101_111_001: wdata <= 1'b0;
      9'b101_111_010: wdata <= 1'b0;
      9'b101_111_011: wdata <= 1'b0;
      9'b101_111_100: wdata <= 1'b0;
      9'b101_111_101: wdata <= 1'b0;
      9'b101_111_110: wdata <= 1'b0;
      9'b101_111_111: wdata <= 1'b0;
      9'b110_000_000: wdata <= 1'b0;
      9'b110_000_001: wdata <= 1'b1;
      9'b110_000_010: wdata <= 1'b1;
      9'b110_000_011: wdata <= 1'b0;
      9'b110_000_100: wdata <= 1'b1;
      9'b110_000_101: wdata <= 1'b0;
      9'b110_000_110: wdata <= 1'b0;
      9'b110_000_111: wdata <= 1'b0;
      9'b110_001_000: wdata <= 1'b1;
      9'b110_001_001: wdata <= 1'b0;
      9'b110_001_010: wdata <= 1'b0;
      9'b110_001_011: wdata <= 1'b0;
      9'b110_001_100: wdata <= 1'b0;
      9'b110_001_101: wdata <= 1'b0;
      9'b110_001_110: wdata <= 1'b0;
      9'b110_001_111: wdata <= 1'b0;
      9'b110_010_000: wdata <= 1'b1;
      9'b110_010_001: wdata <= 1'b1;
      9'b110_010_010: wdata <= 1'b1;
      9'b110_010_011: wdata <= 1'b0;
      9'b110_010_100: wdata <= 1'b1;
      9'b110_010_101: wdata <= 1'b0;
      9'b110_010_110: wdata <= 1'b0;
      9'b110_010_111: wdata <= 1'b0;
      9'b110_011_000: wdata <= 1'b1;
      9'b110_011_001: wdata <= 1'b0;
      9'b110_011_010: wdata <= 1'b0;
      9'b110_011_011: wdata <= 1'b0;
      9'b110_011_100: wdata <= 1'b0;
      9'b110_011_101: wdata <= 1'b0;
      9'b110_011_110: wdata <= 1'b0;
      9'b110_011_111: wdata <= 1'b0;
      9'b110_100_000: wdata <= 1'b1;
      9'b110_100_001: wdata <= 1'b0;
      9'b110_100_010: wdata <= 1'b0;
      9'b110_100_011: wdata <= 1'b0;
      9'b110_100_100: wdata <= 1'b0;
      9'b110_100_101: wdata <= 1'b0;
      9'b110_100_110: wdata <= 1'b0;
      9'b110_100_111: wdata <= 1'b0;
      9'b110_101_000: wdata <= 1'b0;
      9'b110_101_001: wdata <= 1'b0;
      9'b110_101_010: wdata <= 1'b0;
      9'b110_101_011: wdata <= 1'b0;
      9'b110_101_100: wdata <= 1'b0;
      9'b110_101_101: wdata <= 1'b0;
      9'b110_101_110: wdata <= 1'b0;
      9'b110_101_111: wdata <= 1'b0;
      9'b110_110_000: wdata <= 1'b1;
      9'b110_110_001: wdata <= 1'b0;
      9'b110_110_010: wdata <= 1'b0;
      9'b110_110_011: wdata <= 1'b0;
      9'b110_110_100: wdata <= 1'b0;
      9'b110_110_101: wdata <= 1'b0;
      9'b110_110_110: wdata <= 1'b0;
      9'b110_110_111: wdata <= 1'b0;
      9'b110_111_000: wdata <= 1'b0;
      9'b110_111_001: wdata <= 1'b0;
      9'b110_111_010: wdata <= 1'b0;
      9'b110_111_011: wdata <= 1'b0;
      9'b110_111_100: wdata <= 1'b0;
      9'b110_111_101: wdata <= 1'b0;
      9'b110_111_110: wdata <= 1'b0;
      9'b110_111_111: wdata <= 1'b0;
      9'b111_000_000: wdata <= 1'b1;
      9'b111_000_001: wdata <= 1'b0;
      9'b111_000_010: wdata <= 1'b0;
      9'b111_000_011: wdata <= 1'b0;
      9'b111_000_100: wdata <= 1'b0;
      9'b111_000_101: wdata <= 1'b0;
      9'b111_000_110: wdata <= 1'b0;
      9'b111_000_111: wdata <= 1'b0;
      9'b111_001_000: wdata <= 1'b0;
      9'b111_001_001: wdata <= 1'b0;
      9'b111_001_010: wdata <= 1'b0;
      9'b111_001_011: wdata <= 1'b0;
      9'b111_001_100: wdata <= 1'b0;
      9'b111_001_101: wdata <= 1'b0;
      9'b111_001_110: wdata <= 1'b0;
      9'b111_001_111: wdata <= 1'b0;
      9'b111_010_000: wdata <= 1'b1;
      9'b111_010_001: wdata <= 1'b0;
      9'b111_010_010: wdata <= 1'b0;
      9'b111_010_011: wdata <= 1'b0;
      9'b111_010_100: wdata <= 1'b0;
      9'b111_010_101: wdata <= 1'b0;
      9'b111_010_110: wdata <= 1'b0;
      9'b111_010_111: wdata <= 1'b0;
      9'b111_011_000: wdata <= 1'b0;
      9'b111_011_001: wdata <= 1'b0;
      9'b111_011_010: wdata <= 1'b0;
      9'b111_011_011: wdata <= 1'b0;
      9'b111_011_100: wdata <= 1'b0;
      9'b111_011_101: wdata <= 1'b0;
      9'b111_011_110: wdata <= 1'b0;
      9'b111_011_111: wdata <= 1'b0;
      9'b111_100_000: wdata <= 1'b0;
      9'b111_100_001: wdata <= 1'b0;
      9'b111_100_010: wdata <= 1'b0;
      9'b111_100_011: wdata <= 1'b0;
      9'b111_100_100: wdata <= 1'b0;
      9'b111_100_101: wdata <= 1'b0;
      9'b111_100_110: wdata <= 1'b0;
      9'b111_100_111: wdata <= 1'b0;
      9'b111_101_000: wdata <= 1'b0;
      9'b111_101_001: wdata <= 1'b0;
      9'b111_101_010: wdata <= 1'b0;
      9'b111_101_011: wdata <= 1'b0;
      9'b111_101_100: wdata <= 1'b0;
      9'b111_101_101: wdata <= 1'b0;
      9'b111_101_110: wdata <= 1'b0;
      9'b111_101_111: wdata <= 1'b0;
      9'b111_110_000: wdata <= 1'b0;
      9'b111_110_001: wdata <= 1'b0;
      9'b111_110_010: wdata <= 1'b0;
      9'b111_110_011: wdata <= 1'b0;
      9'b111_110_100: wdata <= 1'b0;
      9'b111_110_101: wdata <= 1'b0;
      9'b111_110_110: wdata <= 1'b0;
      9'b111_110_111: wdata <= 1'b0;
      9'b111_111_000: wdata <= 1'b0;
      9'b111_111_001: wdata <= 1'b0;
      9'b111_111_010: wdata <= 1'b0;
      9'b111_111_011: wdata <= 1'b0;
      9'b111_111_100: wdata <= 1'b0;
      9'b111_111_101: wdata <= 1'b0;
      9'b111_111_110: wdata <= 1'b0;
      9'b111_111_111: wdata <= 1'b0;
    endcase
  end // always @ (posedge clk)

endmodule // top
